
configuration topconstruct of top is
  for behave
    for  U1 : cpu use entity work.cpu(EPF10K10TC144_a3);
    end for;
  end for;
end topconstruct;

